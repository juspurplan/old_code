5�d d        d    �� 
 CDflipflop%  i���i  ���                       ��  Cpin%  +���3  +���0 0 CLK  9���        �%  C���3  C���1 1 D1  Q���        �G  i���G  [���1 1 SET';  w���        �G  ���G  ���1 1 RESET'2  ���         �i  C���[  C���0 0 Q1f  Q���        �i  +���[  +���1 1 Q1'f  9���        �$  ����h  7���                       �$  ]���2  ]���0 0 CLK  k���        �$  u���2  u���0 0 D2  ����        �F  ����F  ����1 1 SET':  ����        �F  7���F  E���1 1 RESET'1  7���         �h  u���Z  u���0 0 Q2h  ����        �h  ]���Z  ]���1 1 Q2'h  k���        �3  ����w  E���                       �3  k���A  k���0 0 CLK  y���        �3  ����A  ����0 0 D3#  ����        �U  ����U  ����1 1 SET'I  ����        �U  E���U  S���1 1 RESET'@  E���         �w  ����i  ����0 0 Q3v  ����        �w  k���i  k���1 1 Q3'v  y���        ��  Cswitch&   z���V   n���V   ����n   p��� X     �&   z���4   z���1 1                  �&   n���4   n���0 0                   �V   t���H   t���0 1 XV   ����        �-   `���]   T���]   h����   V��� CLK     �-   `���;   `���1 Z                  �-   T���;   T���0 Z                   �]   Z���O   Z���0 1 CLK]   h���        �0   i���`   ]���`   q����   _��� RESET     �0   i���>   i���1 Z                  �0   ]���>   ]���0 Z                   �`   c���R   c���0 0 RESET`   q���        �� 	 Cinverterl   ^����   :���                       �l   L���z   L���0 0                   ��   L����   L���1 1 X'�   Z���        %��   s����   O���                       ��   a����   a���0 0                   ��   a����   a���1 1 RESET'�   o���        ��  Cor2@  �����  k���                       �@  ����S  ����1 1 X'7  ����        �@  w���S  w���0 0                   ��  }���u  }���1 1 D1�  ����        ��  Cand3�  s���  O���                       ��  m����  m���0 0 Q1�  {���        ��  a����  a���0 0 Q2�  o���        ��  U����  U���1 1 Q3'�  c���         �  a����  a���0 0                  ��  Cor3=  ~����  Z���                       �=  x���P  x���0 0 X6  ����        �=  l���Q  l���0 0 Q1-  z���        �=  `���P  `���0 0 Q2-  n���         ��  l���r  l���0 0 D2�  z���        ��  Cand2�  ����   ����                       ��  �����  ����0 0 X�  ����        ��  �����  ����1 1 Q2'�  ����         �  ����  ����0 0                  =��  T���  0���                       ��  H����  H���1 1 Q1'�  V���        ��  <����  <���0 0 Q2�  J���         �  B���  B���0 0                  ,�<  �����  b���                       �<  z���O  z���0 0                  �<  n���O  n���0 0                   �  t���q  t���0 0 D3  ����        ��  Cand42  ����v  j���                       �2  ����@  ����1 1 X')  ����        �2  ����@  ����1 1 Q1'   ����        �2  v���@  v���0 0 Q2"  ����        �2  j���@  j���1 1 Q3'   x���         �u  |���g  |���0 0 Zu  ����        �0   0���`   $���`   8����   &��� SET     �0   0���>   0���1 Z                  �0   $���>   $���0 1                   �`   *���R   *���0 0 SET`   8���        %��   B����   ���                       ��   0����   0���0 0                   ��   0����   0���1 1 SET'�   >���         ��  Cnet0  ��  Csegmentl   L���l   t���Z�V   t���l   t���Z�V   t���V   t���Z�l   L���l   L��� ' 9 ?   X�0  Z��   a����   c���Z�`   c����   c���Z�`   c���`   c���Z��   a����   a��� *  $ X�1        + X�1    . L  ( X�0    3 :   X�0    4 ; D N   X�1    5 O   X�0  Z�@  w���@  a���Z�  a���@  a���Z�  a���  a���Z�@  w���@  w��� /  6 X�0  Z�<  z���<  ����Z�  ����<  ����Z�  ����  ����Z�<  z���<  z��� G  A X�0  Z�<  n���<  B���Z�  B���<  B���Z�  B���  B���Z�<  n���<  n��� H  E X�1    @   X�1    C M  	 X�1      0 X�0      < X�0      I X�0          X�0  Z��   0����   *���Z�`   *����   *���Z�`   *���`   *���Z��   0����   0��� V  T X�1        W   ajt2459