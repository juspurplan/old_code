library verilog;
use verilog.vl_types.all;
entity Complete_MIPS is
    port(
        CLK             : in     vl_logic;
        RST             : in     vl_logic
    );
end Complete_MIPS;
