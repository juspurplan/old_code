5�� �        d   	 ��  Cand3y  ����  ]���                       ��  Cpiny  �����  ����1 1                  �y  �����  ����0 0                  �y  i����  i���0 0                   ��  �����  ����0 0                  ��  Cand2Y  E����  ����                       �Y  -���u  -���0 0                  �Y  ���u  ���1 1                   ��  !����  !���0 0                  ��  Cor2�  ����{  ����                       ��  ����  ����0 0                  ��  ����  ����0 0                   �y  ����]  ����0 0                  ��  Cswitch#   �����   �����   ����   ���� D     �#   ����?   ����1                    �#   ����?   ����0                     ��   ����g   ����1 0 D�   ���        �   ����w   ����1   ����g   ���� C     �   ����3   ����1                    �   ����3   ����0                     �w   ����[   ����0 0 C1   ����        �   ����o   ����)   ����]   ���� A     �   ����+   ����1                    �   ����+   ����0                     �o   ����S   ����0 0 A)   ����        �   =���}   %���7   a���k   =��� B     �   =���9   =���1                    �   %���9   %���0                     �}   1���a   1���0 0 B7   a���        �� 	 Cinverter  �����  ����                       �  ����)  ����0 0                   ��  ����m  ����1 1                  #��  -����  ����                       ��  	����  	���0 0                   ��  	����  	���1 1                   ��  Cnet0  ��  Csegment�  �����  ����,��  �����  ����,��  �����  ����,��  �����  ����    *�0  ,��  �����  ����,��  -����  ����,��  �����  ����,��  '����  -���,��  -����  -���,��  !����  -���,��  !����  !���    *�0  ,�  ����  ����,��   ����  ����,�o   ����o   ����,�  ����  ����,�o   �����   ����,��   �����   -���,�Y  -����   -���,�Y  -���Y  -��� % 
   *�1  ,�y  ����y  ����,��  ����y  ����,��  �����  ����,�y  ����y  ����   & *�0 
 ,�S  1����  1���,��  o����  1���,�}   1���}   1���,��  o���y  o���,�y  ����y  o���,�y  ����y  ����,�}   1���S  1���,�S  1���S  	���,��  	���S  	���,��  	����  	���  (  " *�0  ,�y  i���y  ����,�y  i���y  i���,�y  ����w   ����,�w   ����w   ����,�w   ����w   ����    *�1  ,�Y  ���Y  	���,��  	���Y  	���,��  	����  	���,�Y  ���Y  ���   )   ajt2459