5�d d        d    �� 
 CDflipflop%  i���i  ���                       ��  Cpin%  +���3  +���0 0 clk  9���        �%  C���3  C���1 1 D1  Q���        �G  i���G  [���1 1                  �G  ���G  ���0 0 rst@  ���         �i  C���[  C���0 0 Q1f  Q���        �i  +���[  +���1 1 Q1'f  9���        �$  ����h  7���                       �$  ]���2  ]���0 0 clk  k���        �$  u���2  u���0 0 D2  ����        �F  ����F  ����1 1                  �F  7���F  E���0 0 rst?  7���         �h  u���Z  u���0 0 Q2h  ����        �h  ]���Z  ]���1 1 Q2'h  k���        �3  ����w  E���                       �3  k���A  k���0 0 clk$  y���        �3  ����A  ����0 0 D3#  ����        �U  ����U  ����1 1                  �U  E���U  S���0 0 rstN  E���         �w  ����i  ����0 0 Q3v  ����        �w  k���i  k���1 1 Q3'v  y���        ��  Cswitch&   z���V   n���V   ����n   p��� X     �&   z���4   z���1 1                  �&   n���4   n���0 0                   �V   t���H   t���0 0 XV   ����        �-   `���]   T���]   h���~   V��� clk     �-   `���;   `���1 Z                  �-   T���;   T���0 Z                   �]   Z���O   Z���0 0 clk]   h���        �0   i���`   ]���`   q����   _��� rst     �0   i���>   i���1 Z                  �0   ]���>   ]���0 Z                   �`   c���R   c���0 0 rst`   q���        �� 	 Cinverterl   ^����   :���                       �l   L���z   L���0 0                   ��   L����   L���1 1 X'�   Z���        ��  Cor2@  �����  k���                       �@  ����S  ����1 1 X'7  ����        �@  w���S  w���0 0                   ��  }���u  }���1 1 D1�  ����        ��  Cand3�  s���  O���                       ��  m����  m���0 0 Q1�  {���        ��  a����  a���0 0 Q2�  o���        ��  U����  U���1 1 Q3'�  c���         �  a����  a���0 0                  ��  Cor3=  ~����  Z���                       �=  x���P  x���0 0 X6  ����        �=  l���Q  l���0 0 Q1-  z���        �=  `���P  `���0 0 Q2-  n���         ��  l���r  l���0 0 D2�  z���        ��  Cand2�  ����   ����                       ��  �����  ����0 0 X�  ����        ��  �����  ����1 1 Q2'�  ����         �  ����  ����0 0                  :��  T���  0���                       ��  H����  H���1 1 Q1'�  V���        ��  <����  <���0 0 Q2�  J���         �  B���  B���0 0                  )�<  �����  b���                       �<  z���O  z���0 0                  �<  n���O  n���0 0                   �  t���q  t���0 0 D3  ����        ��  Cand42  ����v  j���                       �2  ����@  ����1 1 X')  ����        �2  ����@  ����1 1 Q1'   ����        �2  v���@  v���0 0 Q2"  ����        �2  j���@  j���1 1 Q3'   x���         �u  |���g  |���0 0 Zu  ����        ��  Cprobel  �����  |���                        �v  |���v  ����0 0                    N�_  d���s  D���                        �i  D���i  R���0 0                    N�\  ����p  u���                        �f  u���f  ����0 0                    N�j  ����~  ����                        �t  ����t  ����0 0                    ��  CplusV�  �����  ����                          ��  �����  ����1 1                   ��  Cnet0  ��  Csegmentl   L���l   t���\�V   t���l   t���\�V   t���V   t���\�l   L���l   L��� ' 6 <   Z�1      - Z�0  \�i  D���i  C���\�i  D���i  D���\�i  C���i  C��� R 0 7   Z�0  \�@  w���@  a���\�  a���@  a���\�  a���  a���\�@  w���@  w��� ,  3 Z�0  \�<  z���<  ����\�  ����<  ����\�  ����  ����\�<  z���<  z��� D  > Z�0  \�<  n���<  B���\�  B���<  B���\�  B���  B���\�<  n���<  n��� E  B Z�1    @ J  	 Z�0      9 Z�0  \�f  u���h  u���\�f  u���f  u���\�h  u���h  u��� T 1 8 A K   Z�1    =   Z�0      F Z�1    2 L   Z�1    + I  ( Z�0  \�v  |���u  |���\�v  |���v  |���\�u  |���u  |��� P  M Z�0  \�w  ����w  ����\�t  ����w  ����\�t  ����t  ����\�w  ����w  ���� V   Z�1  \�U  ����U  ����\�  ����U  ����\��  �����  ����\�U  ����U  ����\��  ����  ����\�  ����  ����\�  ����  ����\�  ����  ����\�  ����  ����\�B  ����B  ����\�F  ����B  ����\�F  ����F  ����\�B  ����  ����\�  ����  ����\�  ����G  ����\�G  i���G  ����\�G  i���G  i���     Y Z�0  \��   a����   c���\�`   c����   c���\�`   c���`   c���     $ Z�0            ajt2459