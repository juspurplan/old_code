5�d d          ��  Cclock/   -���e   ���e   2����    ���2 CLK       ��  Cpine   $���W   $���1 1 CLKe   2���        �� 
 CDflipflop%  i���i  ���                       �%  +���3  +���1 1 CLK  9���        �%  C���3  C���X X D1  Q���        �G  i���G  [���1 1 SET';  w���        �G  ���G  ���1 1 RESET'2  ���         �i  C���[  C���0 0 Q1f  Q���        �i  +���[  +���1 1 Q1'f  9���        �$  ����h  7���                       �$  ]���2  ]���1 1 CLK  k���        �$  u���2  u���X X D2  ����        �F  ����F  ����1 1 SET':  ����        �F  7���F  E���1 1 RESET'1  7���         �h  u���Z  u���0 0 Q2h  ����        �h  ]���Z  ]���1 1 Q2'h  k���        �3  ����w  E���                       �3  k���A  k���1 1 CLK  y���        �3  ����A  ����X X D3#  ����        �U  ����U  ����1 1 SET'I  ����        �U  E���U  S���1 1 RESET'@  E���         �w  ����i  ����0 0 Q3v  ����        �w  k���i  k���1 1 Q3'v  y���        ��  Cswitch0   i���`   ]���`   q����   _��� RESET     �0   i���>   i���1 Z                  �0   ]���>   ]���0 Z                   �`   c���R   c���0 0 RESET`   q���        �� 	 Cinverter�   s����   O���                       ��   a����   a���0 0                   ��   a����   a���1 1 RESET'�   o���        ��  Cor2@  �����  k���                       �@  ����S  ����X X X'7  ����        �@  w���S  w���0 0                   ��  }���u  }���X X D1�  ����        ��  Cand3�  s���  O���                       ��  m����  m���0 0 Q1�  {���        ��  a����  a���0 0 Q2�  o���        ��  U����  U���1 1 Q3'�  c���         �  a����  a���0 0                  ��  Cor3=  ~����  Z���                       �=  x���P  x���Z Z X6  ����        �=  l���Q  l���0 0 Q1-  z���        �=  `���P  `���0 0 Q2-  n���         ��  l���r  l���X X D2�  z���        ��  Cand2�  ����   ����                       ��  �����  ����Z Z X�  ����        ��  �����  ����1 1 Q2'�  ����         �  ����  ����X X                  5��  T���  0���                       ��  H����  H���1 1 Q1'�  V���        ��  <����  <���0 0 Q2�  J���         �  B���  B���0 0                  $�<  �����  b���                       �<  z���O  z���X X                  �<  n���O  n���0 0                   �  t���q  t���X X D3  ����        ��  Cand42  ����v  j���                       �2  ����@  ����X X X')  ����        �2  ����@  ����1 1 Q1'   ����        �2  v���@  v���0 0 Q2"  ����        �2  j���@  j���1 1 Q3'   x���         �u  |���g  |���0 0 Zu  ����        �0   0���`   $���`   8����   &��� SET     �0   0���>   0���1 Z                  �0   $���>   $���0 1                   �`   *���R   *���0 0 SET`   8���         ��   B����   ���                       ��   0����   0���0 0                   ��   0����   0���1 1 SET'�   >���        ��  Cinput_signal9   ���o   ����F   ���^   ��� X       �o   ����a   ����Z Z Xo   
���         ��  Csignal    Z S�   0 S�}   1 S��   0 S�E  1 S��  0 S�  1 S�q  0 S��  0 S�9  1 S��  0 S�  1 S�e  0 S��  0  ��   �����   ����                       ��   �����   ����Z Z                   ��   �����   ����X X X'�   ����        ��  Cprobey   ����   �����   .����   ���  X     ��   �����   
���Z Z X�   ����          e�[   C���o   #���h   U����   C���  CLK     �e   #���e   1���1 1 CLKY   #���          e�i  ����}  ~���v  �����  ����  Z     �s  ~���s  ����0 0 Zp  ~���          e�]  e���q  E���j  w����  e���  Q1     �g  E���g  S���0 0 Q1_  E���          e�]  ����q  u���j  �����  ����  Q2     �g  u���g  ����0 0 Q2_  u���          e�i  ����}  ����v  �����  ����  Q3     �s  ����s  ����0 0 Q3k  ����           ��  CnetZ  ��  Csegment�   �����   ����t��   �����   ����t�o   ����o   ����t��   �����   ����t�o   �����   ����t��   �����   ���� c g 1 7  R r�0  t��   a����   c���t�`   c����   c���t�`   c���`   c���t��   a����   a��� "   r�X      ( r�1    	    O r�0  t�i  C���i  E���t�g  E���i  E���t�g  E���g  E���t�i  C���i  C��� m + 2   r�0  t�g  u���h  u���t�g  u���g  u���t�h  u���h  u��� o , 3 < F   r�1    
    # r�0  t�@  w���@  a���t�  a���@  a���t�  a���  a���t�@  w���@  w��� '  . r�X  t�<  z���<  ����t�  ����<  ����t�  ����  ����t�<  z���<  z��� ?  9 r�0  t�<  n���<  B���t�  B���<  B���t�  B���  B���t�<  n���<  n��� @  = r�1    ; E   r�X      4 r�1    8   r�X      A r�1    - G   r�1  t�e   #���e   $���t�e   #���e   #���t�e   $���e   $��� i      r�0  t��   0����   *���t�`   *����   *���t�`   *���`   *���t��   0����   0��� N  L r�X    & D  d r�Z       r�0  t�u  |���u  ~���t�s  ~���u  ~���t�s  ~���s  ~���t�u  |���u  |��� k  H r�0  t�w  ����w  ����t�s  ����w  ����t�s  ����s  ����t�w  ����w  ���� q     ajt2459