library verilog;
use verilog.vl_types.all;
entity sorter_testbench is
end sorter_testbench;
