5�d d      �	   ��  Cclock2   ���h   ���?   0���j   ���2 CLK       ��  Cpinh   ���Z   ���1 1 CLKh   #���        �� 
 CDflipflop%  i���i  ���                       �%  +���3  +���1 1 CLK  9���        �%  C���3  C���0 0 D1  Q���        �G  i���G  [���1 1 SET';  w���        �G  ���G  ���1 1 RESET'2  ���         �i  C���[  C���0 0 Q1f  Q���        �i  +���[  +���1 1 Q1'f  9���        �$  ����h  7���                       �$  ]���2  ]���1 1 CLK  k���        �$  u���2  u���1 1 D2  ����        �F  ����F  ����1 1 SET':  ����        �F  7���F  E���1 1 RESET'1  7���         �h  u���Z  u���0 0 Q2h  ����        �h  ]���Z  ]���1 1 Q2'h  k���        �3  ����w  E���                       �3  k���A  k���1 1 CLK  y���        �3  ����A  ����1 1 D3#  ����        �U  ����U  ����1 1 SET'I  ����        �U  E���U  S���1 1 RESET'@  E���         �w  ����i  ����0 0 Q3v  ����        �w  k���i  k���1 1 Q3'v  y���        ��  Cor2@  �����  k���                       �@  ����S  ����0 0 X'7  ����        �@  w���S  w���0 0                   ��  }���u  }���0 0 D1�  ����        ��  Cand3�  s���  O���                       ��  m����  m���0 0 Q1�  {���        ��  a����  a���0 0 Q2�  o���        ��  U����  U���1 1 Q3'�  c���         �  a����  a���0 0                  ��  Cor3=  ~����  Z���                       �=  x���P  x���1 1 X6  ����        �=  l���Q  l���0 0 Q1-  z���        �=  `���P  `���0 0 Q2-  n���         ��  l���r  l���1 1 D2�  z���        ��  Cand2�  ����   ����                       ��  �����  ����1 1 X�  ����        ��  �����  ����1 1 Q2'�  ����         �  ����  ����1 1                  ,��  T���  0���                       ��  H����  H���1 1 Q1'�  V���        ��  <����  <���0 0 Q2�  J���         �  B���  B���0 0                  �<  �����  b���                       �<  z���O  z���1 1                  �<  n���O  n���0 0                   �  t���q  t���1 1 D3  ����        ��  Cand42  ����v  j���                       �2  ����@  ����0 0 X')  ����        �2  ����@  ����1 1 Q1'   ����        �2  v���@  v���0 0 Q2"  ����        �2  j���@  j���1 1 Q3'   x���         �u  |���g  |���0 0 Zu  ����        ��  Cswitch0   0���`   $���`   8����   &��� SET     �0   0���>   0���1 Z                  �0   $���>   $���0 1                   �`   *���R   *���0 0 SET`   8���        �� 	 Cinverter�   B����   ���                       ��   0����   0���0 0                   ��   0����   0���1 1 SET'�   >���        E��   �����   ����                       ��   �����   ����1 1 X�   ����         ��   �����   ����0 0 X'�   ����        ��  Cprobei  ����}  ~���v  �����  ����  Z     �s  ~���s  ����0 0 Zp  ~���          L�]  e���q  E���j  w����  e���  Q1     �g  E���g  S���0 0 Q1_  E���          L�]  ����q  u���j  �����  ����  Q2     �g  u���g  ����0 0 Q2_  u���          L�i  ����}  ����v  �����  ����  Q3     �s  ����s  ����0 0 Q3k  ����          ��  Cchecker�   ����  _���                       ��   �����   ����0 0 Z�   ����        ��   _����   m���1 1 CLK�   _���         ��   �����   ����1 1 RESET'�   ����        �  ����  ����1 1 X  ����        101011101001R010101001010000100000100X000010100000 ��  Cnet1  ��  Csegment�   �����   ����]��   �����   ����]��   �����   ����]�o   �����   ���� ( . J  Z [�1    
    Y [�0     ;  K [�0  ]�i  C���i  E���]�g  E���i  E���]�g  E���g  E���]�i  C���i  C��� " ) P   [�0  ]�g  u���h  u���]�g  u���g  u���]�h  u���h  u��� # * 3 = R   [�1    $ >   [�0  ]�@  w���@  a���]�  a���@  a���]�  a���  a���]�@  w���@  w���   % [�1  ]�<  z���<  ����]�  ����<  ����]�  ����  ����]�<  z���<  z��� 6  0 [�0  ]�<  n���<  B���]�  B���<  B���]�  B���  B���]�<  n���<  n��� 7  4 [�1    /   [�1    2 <   [�0       [�1      + [�1      8 [�1       X   [�0  ]��   0����   *���]�`   *����   *���]�`   *���`   *���]��   0����   0��� G  D [�1     	   H [�Z       [�0  ]�u  |���u  ~���]�s  ~���u  ~���]�s  ~���s  ~���]�u  |���u  |��� N W  ? [�0  ]�w  ����w  ����]�s  ����w  ����]�s  ����s  ����]�w  ����w  ���� T     ajt2459