5�d d        d    ��  Cswitch:   ����j   ����G   ����`   ���� A     ��  Cpin:   ����H   ����1 ��                 �:   ����H   ����0                     �j   ����\   ����1 0 Aj   ����        �D   ����t   ����Q   ���j   ���� B     �D   ����R   ����1 ��                 �D   ����R   ����0 ��                  �t   ����f   ����0 1 Bt   ���        �P   ����   ���]   )���w   ��� C     �P   ���^   ���1 ��                 �P   ���^   ���0 ��                  ��   ���r   ���0 1 C�   ���        �Q   |����   p���^   ����x   |��� D     �Q   |���_   |���1                    �Q   p���_   p���0                     ��   v���s   v���1 1 D�   ����        �H   ����x   ����U   ����n   ���� E     �H   ����V   ����1                    �H   ����V   ����0                     �x   ����j   ����1 1 Ex   ����        �� 	 Cinverter�   �����   m����   �����   ���� A'     ��   ����   ���1 1                   ��   ����   ���0 0                  ��   �����   �����   �����   ���� B'     ��   �����   ����0 0                   ��   �����   ����1 1                  ��   6����   ����   H����   6��� D'     ��   $����   $���1 1                   ��   $����   $���0 0                  ��   f����   B����   x����   f��� E'     ��   T����   T���1 1                   ��   T����   T���0 0                  ��  Cnor3  ����Q  ����  ����O  ���� A+B+C     �  ����  ����1 1                  �  ����  ����0 0                  �  ����  ����0 0                   �P  ����B  ����0 0                  $�	  }���T  Y���  ����R  }��� A+C+E     �	  w���  w���1 1                  �	  k���  k���0 0                  �	  _���  _���1 1                   �S  k���E  k���0 0                  $�  9���R  ���  K���S  9��� A'+C+E     �  3���  3���0 0                  �  '���  '���0 0                  �  ���  ���1 1                   �Q  '���C  '���0 0                  $�  ����Q  ����  ����U  ���� B'+C+E'     �  ����  ����1 1                  �  ����  ����0 0                  �  ����  ����0 0                   �P  ����B  ����0 0                  $�   ����K  |���  ����I  ���� A+B+D     �   ����  ����1 1                  �   ����  ����0 0                  �   ����  ����1 1                   �J  ����<  ����0 0                  $�  =���R  ���  O���Q  =��� C+D+E     �  7���  7���0 0                  �  +���  +���1 1                  �  ���  ���1 1                   �Q  +���C  +���0 0                  $�  ����P  ����  ����T  ���� A'+B'+D     �  ����  ����0 0                  �  ����  ����1 1                  �  ����  ����1 1                   �O  ����A  ����0 0                  $�  /���P  ���  A���M  /��� A+B+E     �  )���  )���1 1                  �  ���  ���0 0                  �  ���  ���1 1                   �O  ���A  ���0 0                  $�  ����L  ����  ����N  ���� A'+C+D     �  ����  ����0 0                  �  ����  ����0 0                  �  ����  ����1 1                   �K  ����=  ����0 0                  $�
  p���U  L���  ����S  p��� A+D+E     �
  j���  j���1 1                  �
  ^���  ^���1 1                  �
  R���  R���1 1                   �T  ^���F  ^���0 0                  ��  Cnor4  ����V  i���  ����o  ���� 
B'+C+D'+E'     �  ����  ����1 1                  �  ����  ����0 0                  �  u���  u���0 0                  �  i���  i���0 0                   �U  {���G  {���0 0                  W�`  �����  s���m  �����  ���� W     �`  ����n  ����0 0                  �`  ����s  ����0 0                  �`  ���s  ���0 0                  �`  s���n  s���0 0                   ��  �����  ����1 1                  W�5  �����  ����B  ����Z  ���� Z     �5  ����C  ����0 0                  �5  ����H  ����0 0                  �5  ����H  ����0 0                  �5  ����C  ����0 0                   �  ����q  ����1 1                  ��  Cnor5$  ����o  ����.  ����F  ���� X     �$  ����2  ����0 0                  �$  ����7  ����0 0                  �$  ����8  ����0 0                  �$  ����7  ����0 0                  �$  ����2  ����0 0                   �n  ����`  ����1 1                  j�  ����d  ����&  ����?  ���� Y     �  ����'  ����0 0                  �  ����,  ����0 0                  �  ����-  ����0 0                  �  ����,  ����0 0                  �  ����'  ����0 0                   �c  ����U  ����1 1                  ��  Cnor2	  ���T  ����  $���F  ��� A'+B'     �	  ���  ���0 0                  �	  ����  ����1 1                   �S   ���E   ���0 0                  y�  ����Z  ����  ����H  ���� C+D     �  ����"  ����0 0                  �  ����"  ����1 1                   �Y  ����K  ����0 0                  y�  {���]  W���  ����J  {��� C+E     �  o���%  o���0 0                  �  c���%  c���1 1                   �\  i���N  i���0 0                  y�  <���_  ���!  N���K  <��� A+B     �  0���'  0���1 1                  �  $���'  $���0 0                   �^  *���P  *���0 0                   ��  Cnet1  ��  Csegment�   ����   ������j   �����   ������j   ����j   �������   ����   �����  �����   ������  0���  �����  ����  ������  ����  ������  ����  ������  w���	  w�����  ����  w�����	  w���	  w�����  ����   ������  w���  ������   ����   ������  )���  )�����  )���  )�����  j���
  j�����  )���  j�����
  j���
  j�����  0���  0�����  j���  0�����  0���  0�����  )���  ����  & + : I S �   ��0  ���   �����   �������   �����   �������   �����   �������   �����   �������   �����   ������t   �����   ������t   ����t   ������<  �����   ������<  $���<  �����<  ����<  ������<  ����  ������<  ����<  ������  ����  ������<  ����   ������<  ����<  ������   ����   ������<  ���  �����<  ����<  �����  ���  �����<  $���  $�����  $���  $�����<  $���<  ���  ' ; J �  
 ��1  ���   $����   v������   v����   v������   v����   v������   $����   $������   v����   {������  {����   {������  �����  ������  �����  �������  ����   �������  +����  ������   ����   �������  +���  +������  �����  +�����  +���  +������  ����  �������  {����  ������  ����  �������  ^���
  ^������  �����  ^�����
  ^���
  ^������  ����  �������  ^����  ������  ����  �������  ����  �������  {����  ������  ����  ����  < @ F T � P   ��1  ���   T����   ������x   �����   ������x   ����x   �������   T����   T������   �����  �������  ����  �������  _���	  _������  �����  _�����	  _���	  _������  ���  ������  _����  �����  ���  ������  ���  �����  ���  ������  ���  ������  ����  �����  ���  ������  F����  �������  c����  F�����
  F����  F�����
  R���
  F�����
  R���
  R������  c���  c������  �����  c�����  c���  c������  ����  ��� " - 2 A K U �   ��Z       ��Z       ��Z       ��Z       ��0  ���   ���&  �����&  3���&  ������   ����   �����&  ���&  ������&  3���  3�����&  ����&  3�����  3���  3�����&  ����  ������&  ����&  ������  ����  ������&  ����  ������&  ���&  ������  ����  ������&  ���	  �����&  ���&  �����	  ���	  ��� 0 D N {   ��0   ���   ���o  �����o  ����o  ������   ����   �����o  ����o  ������j  ����o  ������o  ����  ������o  k���o  ������  ����  ������o  k���	  k�����o  '���o  k�����	  k���	  k�����o  '���  '�����o  ����o  '�����  '���  '�����o  ����  ������o  7���o  ������  ����  ������o  7���  7�����o  ���o  7�����  7���  7�����o  ����  ������  ����  ������o  ����  ������o  o���o  ������  ����  ������o  o���  o�����o  ���o  o�����  o���  o�����o  ����o  ������o  ����  ������o  ����o  ������  ����  ����	 ( , 1 6 ? Z  � O   ��0  ���   $����  $������  ����  $������   $����   $������  u����  �������  u���  u������  $����  u�����  u���  u��� [    ��0 
 ���   T����  T������  �����  T������   T����   T������  i����  T������  i���  i������  �����  i�����  i���  i������  ����  �������  �����  ������  ����  ���� \ 7  # ��0  ��P  ����P  ������`  ����`  ������P  ����P  ������`  ����P  ���� _  ) ��0  ��S  ����S  k�����`  ����`  ������S  k���S  k�����`  ����S  ���� `  . ��0  ��Q  '���Q  '�����Q  '���Q  %�����Q  '���Q  '�����Q  ,���Q  '������  �����  ,�����$  ����$  �������  ,���Q  ,�����$  �����  ���� l  3 ��0  ��5  ����5  �������  �����  i�����\  i����  i�����\  i���\  i�����5  �����  ���� f  � ��0  ��P  ����P  ������$  ����$  ������P  ����P  ������$  ����P  ���� m  8 ��0  ���  �����  ������  ����  �������  ����U  ������U  {���U  ������U  {���U  {�����  �����  ���� t  ] ��0  ���  �����  �����  ����  �������  ���O  �����O  ���O  �����O  ���O  �����  �����  ���� u  L ��0  ���  �����  ������  ����  �������  ����K  ������K  ����K  ������K  ����K  ������  �����  ���� v  Q ��0  ��  ����  b�����  ����  ������  _���T  _�����T  ^���T  _�����T  ^���T  ^�����  _���  b������  b���  b������  �����  b�����5  ����5  ������  ����  ������5  �����  ���� w h  V ��1  ��	  ����	  ������V  ����	  ������V  ����V  ������   ����V  ������V  ����V  �������   �����   ������V  ����V  ������V  ����V  ������  ����V  ������  ����  ������  ����  ������V  ����  ������  ����  ������V  ����V  ������V  ����  ������V  ����V  ������  ����  ���� | 5 E Y   ��0  ��`  s���`  s�����y  s���y  ������Y  ����y  ������Y  ����Y  ������`  s���y  s��� b  � ��0  ��`  ���`  �����a  ���a   �����S   ���a   �����S   ���S   ������   ���a   �����$  ����$  �������  �����   ������   ����   �����5  ����5  �������  �����   �����`  ���a  �����$  �����  ������5  �����  ���� a p e  } ��0  ��$  ����$  �������  �����  �������  �����  �������  ����J  ������J  ����J  ������$  �����  ���� n  = ��0 	 ��$  ����$  �������  �����  8������  -����  8������  -����  .�����Q  .����  .�����a  .���Q  .�����Q  +���Q  .�����Q  +���Q  +�����$  �����  ���� o  B ��Z  ���  �����  �������  �����  ����    ��0  ��O  ����O  ������O  �����  �������  �����  �������  �����  ������  ����  ������  �����  ���� s  G ��Z       ��0  ��5  ����5  �������  �����  *�����^  *����  *�����^  *���^  *�����5  �����  ���� g  �   ajt2459