5�d d        d    �� 
 CDflipflop%  i���i  ���                       ��  Cpin%  +���3  +���0 0 CLK  9���        �%  C���3  C���1 1 D1  Q���        �G  i���G  [���1 1 SET';  w���        �G  ���G  ���1 1 RESET'2  ���         �i  C���[  C���0 0 Q1f  Q���        �i  +���[  +���1 1 Q1'f  9���        �$  ����h  7���                       �$  ]���2  ]���0 0 CLK  k���        �$  u���2  u���0 0 D2  ����        �F  ����F  ����1 1 SET':  ����        �F  7���F  E���1 1 RESET'1  7���         �h  u���Z  u���0 0 Q2h  ����        �h  ]���Z  ]���1 1 Q2'h  k���        �3  ����w  E���                       �3  k���A  k���0 0 CLK  y���        �3  ����A  ����0 0 D3#  ����        �U  ����U  ����1 1 SET'I  ����        �U  E���U  S���1 1 RESET'@  E���         �w  ����i  ����0 0 Q3v  ����        �w  k���i  k���1 1 Q3'v  y���        ��  Cswitch&   z���V   n���V   ����n   p��� X     �&   z���4   z���1 1                  �&   n���4   n���0 0                   �V   t���H   t���0 0 XV   ����        �-   `���]   T���]   h����   V��� CLK     �-   `���;   `���1 Z                  �-   T���;   T���0 Z                   �]   Z���O   Z���0 0 CLK]   h���        �0   i���`   ]���`   q����   _��� RESET     �0   i���>   i���1 Z                  �0   ]���>   ]���0 Z                   �`   c���R   c���0 0 RESET`   q���        �� 	 Cinverterl   ^����   :���                       �l   L���z   L���0 0                   ��   L����   L���1 1 X'�   Z���        %��   s����   O���                       ��   a����   a���0 0                   ��   a����   a���1 1 RESET'�   o���        ��  Cor2@  �����  k���                       �@  ����S  ����1 1 X'7  ����        �@  w���S  w���0 0                   ��  }���u  }���1 1 D1�  ����        ��  Cand3�  s���  O���                       ��  m����  m���0 0 Q1�  {���        ��  a����  a���0 0 Q2�  o���        ��  U����  U���1 1 Q3'�  c���         �  a����  a���0 0                  ��  Cor3=  ~����  Z���                       �=  x���P  x���0 0 X6  ����        �=  l���Q  l���0 0 Q1-  z���        �=  `���P  `���0 0 Q2-  n���         ��  l���r  l���0 0 D2�  z���        ��  Cand2�  ����   ����                       ��  �����  ����0 0 X�  ����        ��  �����  ����1 1 Q2'�  ����         �  ����  ����0 0                  =��  T���  0���                       ��  H����  H���1 1 Q1'�  V���        ��  <����  <���0 0 Q2�  J���         �  B���  B���0 0                  ,�<  �����  b���                       �<  z���O  z���0 0                  �<  n���O  n���0 0                   �  t���q  t���0 0 D3  ����        ��  Cand42  ����v  j���                       �2  ����@  ����1 1 X')  ����        �2  ����@  ����1 1 Q1'   ����        �2  v���@  v���0 0 Q2"  ����        �2  j���@  j���1 1 Q3'   x���         �u  |���g  |���0 0 Zu  ����        �0   0���`   $���`   8����   &��� SET     �0   0���>   0���1 Z                  �0   $���>   $���0 1                   �`   *���R   *���0 0 SET`   8���        %��   B����   ���                       ��   0����   0���0 0                   ��   0����   0���1 1 SET'�   >���        ��  Cprobel  �����  |���                        �v  |���v  ����0 0                    X�_  d���s  D���                        �i  D���i  R���0 0                    X�\  ����p  u���                        �f  u���f  ����0 0                    X�j  ����~  ����                        �t  ����t  ����0 0                     ��  Cnet0  ��  Csegmentl   L���l   t���c�V   t���l   t���c�V   t���V   t���c�l   L���l   L��� ' 9 ?   a�0  c��   a����   c���c�`   c����   c���c�`   c���`   c���c��   a����   a��� *  $ a�0          a�1      0 a�1        W a�1        + a�0  c�i  D���i  C���c�i  D���i  D���c�i  C���i  C��� 3 : \   a�0  c�@  w���@  a���c�  a���@  a���c�  a���  a���c�@  w���@  w��� /  6 a�0  c�<  z���<  ����c�  ����<  ����c�  ����  ����c�<  z���<  z��� G  A a�0  c�<  n���<  B���c�  B���<  B���c�  B���  B���c�<  n���<  n��� H  E a�1    C M  	 a�0      < a�0  c�f  u���h  u���c�f  u���f  u���c�h  u���h  u��� 4 ; D N ^   a�1    @   a�0      I a�1    5 O   a�0  c��   0����   *���c�`   *����   *���c�`   *���`   *���c��   0����   0��� V  T a�1    . L  ( a�0  c�v  |���u  |���c�v  |���v  |���c�u  |���u  |��� Z  P a�0  c�w  ����w  ����c�t  ����w  ����c�t  ����t  ����c�w  ����w  ���� `     ajt2459