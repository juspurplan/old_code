5�d d        d     ��  Cswitch:   ����j   ����j   �����   ���� A     ��  Cpin:   ����H   ����1 ��                 �:   ����H   ����0                     �j   ����\   ����1 1 Aj   ����        �D   ����t   ����t   ����   ���� B     �D   ����R   ����1 ��                 �D   ����R   ����0 ��                  �t   ����f   ����0 0 Bt   ���        �P   ����   ����   ����   ��� C     �P   ���^   ���1 ��                 �P   ���^   ���0 ��                  ��   ���r   ���0 0 C�   ���        �Q   |����   p����   �����   r��� D     �Q   |���_   |���1                    �Q   p���_   p���0                     ��   v���s   v���1 1 D�   ����        �H   ����x   ����x   �����   ���� E     �H   ����V   ����1                    �H   ����V   ����0                     �x   ����j   ����1 1 Ex   ����        �� 	 Cinverter�   �����   m���                       ��   ����   ���1 1                   ��   ����   ���0 0 A'�   ����        ��   �����   ����                       ��   �����   ����0 0                   ��   �����   ����1 1 B'�   ����        ��   6����   ���                       ��   $����   $���1 1                   ��   $����   $���0 0 D'�   2���        ��   f����   B���                       ��   T����   T���1 1                   ��   T����   T���0 0 E'�   b���        ��  Cnor3  ����Q  ����  ����O  ���� A+B+C     �  ����  ����1 1 A�  ����        �  ����  ����0 0 B�  ����        �  ����  ����0 0 C�  ����         �P  ����B  ����0 0                  $�	  }���T  Y���  ����R  }��� A+C+E     �	  w���  w���1 1 A  ����        �	  k���  k���0 0 C   y���        �	  _���  _���1 1 E  m���         �S  k���E  k���0 0                  $�  9���R  ���  K���S  9��� A'+C+E     �  3���  3���0 0 A'�  A���        �  '���  '���0 0 C�  5���        �  ���  ���1 1 E�  )���         �Q  '���C  '���0 0                  $�  ����Q  ����  ����U  ���� B'+C+E'     �  ����  ����1 1 B'�  ����        �  ����  ����0 0 C�  ����        �  ����  ����0 0 E'�  ����         �P  ����B  ����0 0                  $�   ����K  |���  ����I  ���� A+B+D     �   ����  ����1 1 A�  ����        �   ����  ����0 0 B�  ����        �   ����  ����1 1 D�  ����         �J  ����<  ����0 0                  $�  =���R  ���  O���Q  =��� C+D+E     �  7���  7���0 0 C�  E���        �  +���  +���1 1 D�  9���        �  ���  ���1 1 E�  -���         �Q  +���C  +���0 0                  $�  ����P  ����  ����T  ���� A'+B'+D     �  ����  ����0 0 A'�  ����        �  ����  ����1 1 B'�  ����        �  ����  ����1 1 D�  ����         �O  ����A  ����0 0                  $�  /���P  ���  A���M  /��� A+B+E     �  )���  )���1 1 A�  7���        �  ���  ���0 0 B�  +���        �  ���  ���1 1 E�  ���         �O  ���A  ���0 0                  $�  ����L  ����  ����N  ���� A'+C+D     �  ����  ����0 0 A'�  ����        �  ����  ����0 0 C�  ����        �  ����  ����1 1 D�  ����         �K  ����=  ����0 0                  $�
  p���U  L���  ����S  p��� A+D+E     �
  j���  j���1 1 A  x���        �
  ^���  ^���1 1 D  l���        �
  R���  R���1 1 E  `���         �T  ^���F  ^���0 0                  ��  Cnor4  ����V  i���  ����o  ���� 
B'+C+D'+E'     �  ����  ����1 1 B'  ����        �  ����  ����0 0 C  ����        �  u���  u���0 0 D'   ����        �  i���  i���0 0 E'  w���         �U  {���G  {���0 0                  W�`  �����  s���m  �����  ���� W     �`  ����n  ����0 0                  �`  ����s  ����0 0                  �`  ���s  ���0 0                  �`  s���n  s���0 0                   ��  �����  ����1 1                  W�5  �����  ����B  ����Z  ���� Z     �5  ����C  ����0 0                  �5  ����H  ����0 0                  �5  ����H  ����0 0                  �5  ����C  ����0 0                   �  ����q  ����1 1                  ��  Cnor5$  ����o  ����.  ����F  ���� X     �$  ����2  ����0 0                  �$  ����7  ����0 0                  �$  ����8  ����0 0                  �$  ����7  ����0 0                  �$  ����2  ����0 0                   �n  ����`  ����1 1                  j�  ����d  ����&  ����?  ���� Y     �  ����'  ����0 0                  �  ����,  ����0 0                  �  ����-  ����0 0                  �  ����,  ����0 0                  �  ����'  ����0 0                   �c  ����U  ����1 1                  ��  Cnor2	  ���T  ����  $���F  ��� A'+B'     �	  ���  ���0 0 A'   ���        �	  ����  ����1 1 B'�  ���         �S   ���E   ���0 0                  y�  ����Z  ����  ����H  ���� C+D     �  ����"  ����0 0 C  ����        �  ����"  ����1 1 D  ����         �Y  ����K  ����0 0                  y�  {���]  W���  ����J  {��� C+E     �  o���%  o���0 0 C	  }���        �  c���%  c���1 1 E
  q���         �\  i���N  i���0 0                  y�  <���_  ���!  N���K  <��� A+B     �  0���'  0���1 1 A  >���        �  $���'  $���0 0 B  2���         �^  *���P  *���0 0                  ��  Cprobe�  �����  �����  �����  ����  W     ��  �����  ����1 1 W�  ����          ��a  ����u  ����n  �����  ����  X     �k  ����k  ����1 1 Xh  ����          ��V  ����j  ����c  ����|  ����  Y     �`  ����`  ����1 1 Y]  ����          ��r  �����  ����  �����  ����  Z     �|  ����|  ����1 1 Zy  ����          $ ��  Cnet1  ��  Csegment�   ����   ������   ����   ������j   �����   ������  �����   ������  ����  ������j   ����j   ����  & + : I S �   ��1  ���   $����   v������   v����   v������   v����   v������   $����   $������   v����   {���  < @ F P T �   ��0   	 ( , 1 6 ? O Z  �   ��0    0 D N {   ��1    5 E Y |   ��0    [    ��0  ��P  ����P  ������`  ����`  ������P  ����P  ������`  ����P  ���� _  ) ��0  ��S  ����S  k�����`  ����`  ������S  k���S  k�����`  ����S  ���� `  . ��0  ��Q  '���Q  '�����Q  '���Q  %�����Q  '���Q  '�����Q  ,���Q  '������  �����  ,�����$  ����$  �������  ,���Q  ,�����$  �����  ���� l  3 ��0  ��5  ����5  �������  �����  i�����\  i����  i�����\  i���\  i�����5  �����  ���� f  � ��0  ��P  ����P  ������$  ����$  ������P  ����P  ������$  ����P  ���� m  8 ��0  ���  �����  ������  ����  �������  ����U  ������U  {���U  ������U  {���U  {�����  �����  ���� t  ] ��0  ���  �����  �����  ����  �������  ���O  �����O  ���O  �����O  ���O  �����  �����  ���� u  L ��0  ���  �����  ������  ����  �������  ����K  ������K  ����K  ������K  ����K  ������  �����  ���� v  Q ��0  ��  ����  b�����  ����  ������  _���T  _�����T  ^���T  _�����T  ^���T  ^�����  _���  b������  b���  b������  �����  b�����5  ����5  ������  ����  ������5  �����  ���� w h  V ��0  ��`  s���`  s�����y  s���y  ������Y  ����y  ������Y  ����Y  ������`  s���y  s��� b  � ��0  ��`  ���`  �����a  ���a   �����S   ���a   �����S   ���S   ������   ���a   �����$  ����$  �������  �����   ������   ����   �����5  ����5  �������  �����   �����`  ���a  �����$  �����  ������5  �����  ���� a p e  } ��0  ��$  ����$  �������  �����  �������  �����  �������  ����J  ������J  ����J  ������$  �����  ���� n  = ��0 	 ��$  ����$  �������  �����  8������  -����  8������  -����  .�����Q  .����  .�����a  .���Q  .�����Q  +���Q  .�����Q  +���Q  +�����$  �����  ���� o  B ��Z  ���  �����  �������  �����  ����    ��0  ��O  ����O  ������O  �����  �������  �����  �������  �����  ������  ����  ������  �����  ���� s  G ��0    7 \  # ��0  ��5  ����5  �������  �����  *�����^  *����  *�����^  *���^  *�����5  �����  ���� g  � ��Z  ��j  ����o  ����    ��Z       ��0       ��0       ��0  ���   �����   �������   �����   �������   �����   �������   �����   ������t   �����   ������t   ����t   ����  ' ; J �  
 ��1       ��0       ��0       ��1  ���   T����   T������   T����   ������x   �����   ������x   ����x   ���� " - 2 A K � U   ��1  ���  �����  �������  �����  �������  �����  �������  �����  ���� �  c ��1  ��k  ����n  ������k  ����k  ������n  ����n  ���� �  q ��1  ��`  ����c  ������`  ����`  ������c  ����c  ���� �  x ��1  ��  ����  ������|  ����  ������|  ����|  ������  ����  ���� �  i   ajt2459